//alu parametrizable de n bits. Recibirá dos entradas de n bits y un bus de control