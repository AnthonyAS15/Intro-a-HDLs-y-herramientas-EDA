`timescale 1ns/1ps

module tb_encoder_decoder();

reg [3:0] d;
wire s_a, s_b, s_c, s_d, s_e, s_f, s_g;

seven_segment_display_deco dut(d, s_a, s_b, s_c, s_d, s_e, s_f, s_g);

initial begin

d = 4'b0000; #10;
d = 4'b0001; #10;
d = 4'b0010; #10;
d = 4'b0011; #10;
d = 4'b0100; #10;
d = 4'b0101; #10;
d = 4'b0110; #10;
d = 4'b0111; #10;
d = 4'b1000; #10;
d = 4'b1001; #10;
d = 4'b1010; #10;
d = 4'b1011; #10;
d = 4'b1100; #10;
d = 4'b1101; #10;
d = 4'b1110; #10;
d = 4'b1111; #10;

$finish;

end

endmodule
